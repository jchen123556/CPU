module decoder_6_64(input [5:0] in, [63:0] out);
reg [63:0] out_reg;

always @(*) begin
case (in)
6'h0 : out_reg = 64'h0000000000000001;
6'h1 : out_reg = 64'h0000000000000002;
6'h2 : out_reg = 64'h0000000000000004;
6'h3 : out_reg = 64'h0000000000000008;
6'h4 : out_reg = 64'h0000000000000010;
6'h5 : out_reg = 64'h0000000000000020;
6'h6 : out_reg = 64'h0000000000000040;
6'h7 : out_reg = 64'h0000000000000080;
6'h8 : out_reg = 64'h0000000000000100;
6'h9 : out_reg = 64'h0000000000000200;
6'ha : out_reg = 64'h0000000000000400;
6'hb : out_reg = 64'h0000000000000800;
6'hc : out_reg = 64'h0000000000001000;
6'hd : out_reg = 64'h0000000000002000;
6'he : out_reg = 64'h0000000000004000;
6'hf : out_reg = 64'h0000000000008000;
6'h10 : out_reg = 64'h0000000000010000;
6'h11 : out_reg = 64'h0000000000020000;
6'h12 : out_reg = 64'h0000000000040000;
6'h13 : out_reg = 64'h0000000000080000;
6'h14 : out_reg = 64'h0000000000100000;
6'h15 : out_reg = 64'h0000000000200000;
6'h16 : out_reg = 64'h0000000000400000;
6'h17 : out_reg = 64'h0000000000800000;
6'h18 : out_reg = 64'h0000000001000000;
6'h19 : out_reg = 64'h0000000002000000;
6'h1a : out_reg = 64'h0000000004000000;
6'h1b : out_reg = 64'h0000000008000000;
6'h1c : out_reg = 64'h0000000010000000;
6'h1d : out_reg = 64'h0000000020000000;
6'h1e : out_reg = 64'h0000000040000000;
6'h1f : out_reg = 64'h0000000080000000;
6'h20 : out_reg = 64'h0000000100000000;
6'h21 : out_reg = 64'h0000000200000000;
6'h22 : out_reg = 64'h0000000400000000;
6'h23 : out_reg = 64'h0000000800000000;
6'h24 : out_reg = 64'h0000001000000000;
6'h25 : out_reg = 64'h0000002000000000;
6'h26 : out_reg = 64'h0000004000000000;
6'h27 : out_reg = 64'h0000008000000000;
6'h28 : out_reg = 64'h0000010000000000;
6'h29 : out_reg = 64'h0000020000000000;
6'h2a : out_reg = 64'h0000040000000000;
6'h2b : out_reg = 64'h0000080000000000;
6'h2c : out_reg = 64'h0000100000000000;
6'h2d : out_reg = 64'h0000200000000000;
6'h2e : out_reg = 64'h0000400000000000;
6'h2f : out_reg = 64'h0000800000000000;
6'h30 : out_reg = 64'h0001000000000000;
6'h31 : out_reg = 64'h0002000000000000;
6'h32 : out_reg = 64'h0004000000000000;
6'h33 : out_reg = 64'h0008000000000000;
6'h34 : out_reg = 64'h0010000000000000;
6'h35 : out_reg = 64'h0020000000000000;
6'h36 : out_reg = 64'h0040000000000000;
6'h37 : out_reg = 64'h0080000000000000;
6'h38 : out_reg = 64'h0100000000000000;
6'h39 : out_reg = 64'h0200000000000000;
6'h3a : out_reg = 64'h0400000000000000;
6'h3b : out_reg = 64'h0800000000000000;
6'h3c : out_reg = 64'h1000000000000000;
6'h3d : out_reg = 64'h2000000000000000;
6'h3e : out_reg = 64'h4000000000000000;
6'h3f : out_reg = 64'h8000000000000000;
default : out_reg = 64'h0000000000000000;
endcase
end
assign out = out_reg;
endmodule

module decoder_3_8(input [2:0] in, [7:0] out);
reg [15:0] out_reg;
always @(*) begin
case (in)
3'b000 : out_reg = 8'h01;
3'b001 : out_reg = 8'h02;
3'b010 : out_reg = 8'h04;
3'b011 : out_reg = 8'h08;
3'b100 : out_reg = 8'h10;
3'b101 : out_reg = 8'h20;
3'b110 : out_reg = 8'h40;
3'b111 : out_reg = 8'h80;
default : out_reg = 8'b00;
endcase
end
assign out = out_reg;
endmodule